library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package cl10_fifo_pkg is

end package cl10_fifo_pkg;
