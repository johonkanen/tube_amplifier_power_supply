library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package uart_commands is

    type t_system_states is (eka,toka,kolmas);
    signal st_system_states : t_system_states;


    constant unsigned(15 downto 0) 

end uart_commands;
