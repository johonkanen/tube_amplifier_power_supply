library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package onboard_ad_control_internal_pkg is

end package onboard_ad_control_internal_pkg;
