library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package alu16bit_pkg is

   type t_alu_commands is (nop,add,sub,a_mpy_b,a_div_b,sqrt_a);

end package;
